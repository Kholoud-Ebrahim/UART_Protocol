package param_pkg;
    parameter DWIDTH =6;
    parameter PERIOD = 5;
endpackage :param_pkg