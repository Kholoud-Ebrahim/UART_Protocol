package param_pkg;
    parameter DWIDTH   = 8;
    parameter PWIDTH   = 6; 
    parameter PRESCALE = 8;

    parameter TXPERIOD = 80; // RXPERIOD*PRESCALE
    parameter RXPERIOD = 10; 
endpackage :param_pkg